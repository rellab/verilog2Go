module adder(a, b, q);
input [3:0] a, b;
output [0:3] q;

assign q = 4'b1100;

endmodule